module tdata_acquire;
reg clk_i, reset_n_i, adc_data_rdy_i, syncro_i;
reg [11:0] adc_data_i;
reg adc_data_i_flag;
wire [11:0]	data_o;
wire data_rdy_o;
//????????????? ????????? ???????????? ?????? data_acquire
data_acquire inst(clk_i, reset_n_i, adc_data_req_o, adc_data_rdy_i, adc_data_i, syncro_i, data_o, data_rdy_o);

//adc inst2(clk_i, reset_n_i, adc_data_req_o, adc_data_rdy_i, adc_data_i);
 
 //?????????? ?????? ???????? ??????? 
always#10 clk_i = ~clk_i;
 //?? ?????? ???????... 
initial begin
clk_i = 0; 
reset_n_i = 1; 
adc_data_i = 12'h00;
adc_data_rdy_i = 1'b0; 
syncro_i=1'b0;

//????? ????????? ???????? "50" ?????? ?????? ?????? 
#50 reset_n_i = 0; 
//??? ????? ????? "4" ??????? ?????? ??????
#4 reset_n_i = 1;
//????? ????????????? "50"
 #50; 
//???? ?????? ???????? ??????? ? ????? ????? ??? ?????? ?????? ??????
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-512; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end

//-------------------------------
// ?????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-312; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------
//-------------------------------
// ?????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-157; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------
//-------------------------------
// ????????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-200; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------

//-------------------------------
// ????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-700; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------
//-------------------------------
// ?????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-20; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------


//-------------------------------
// ??????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=-920; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------

//-------------------------------
// ??????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=820; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------

//-------------------------------
// ??????? ?????????
//-------------------------------
@(posedge clk_i)
#20 begin 
syncro_i = 1'b1;
adc_data_rdy_i=0;
end
//?? ?????????? ?????? ??????? ?????? ?????? 
@(posedge clk_i)
#80 begin 
syncro_i = 1'b0;
end

@(negedge adc_data_req_o)
#0 begin
adc_data_i_flag =1;
end

@(posedge clk_i)
#0 begin 
if(adc_data_i_flag) begin #10 begin adc_data_i=1020; end end
end

@(posedge clk_i)
#20 begin 
adc_data_rdy_i=1;
adc_data_i_flag =0;
end
//----------------------------------
end 
//??????????? ????????? ? ?????? ??????? "3400" 
initial begin
#4400 $finish;
end
//??????? ???? VCD ??? ???????????? ??????? ????????
//initial begin $dumpfile("out.vcd");
//$dumpvars(0,test_counter);
//end 
//????????? ?? ?????????? ????????? ??????? 
initial $monitor($stime,, reset_n_i,, clk_i,,, adc_data_req_o);
endmodule